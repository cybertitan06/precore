   module ID_S_5d0f61ec_7e71e69b_E (output reg ID_S_2b616_71_E, input ID_S_2b609_64_E, input clock, input reset); always @(posedge clock) begin if (reset == 1) begin ID_S_2b616_71_E <= 0; end else begin ID_S_2b616_71_E <= ID_S_2b609_64_E; end end endmodule module ID_S_7efb9f9e_394c97fa_E (input [3:0] ID_S_108d5742_7edd6db7_E, output reg [7:0] ID_S_192fd704_45804608_E, input clock); always @(posedge clock) begin case (ID_S_108d5742_7edd6db7_E) 4'b0000: ID_S_192fd704_45804608_E <= 8'b01000000; 4'b0001: ID_S_192fd704_45804608_E <= 8'b01111001; 4'b0010: ID_S_192fd704_45804608_E <= 8'b00100100; 4'b0011: ID_S_192fd704_45804608_E <= 8'b00110000; 4'b0100: ID_S_192fd704_45804608_E <= 8'b00011001; 4'b0101: ID_S_192fd704_45804608_E <= 8'b00010010; 4'b0110: ID_S_192fd704_45804608_E <= 8'b00000010; 4'b0111: ID_S_192fd704_45804608_E <= 8'b01111000; 4'b1000: ID_S_192fd704_45804608_E <= 8'b00000000; 4'b1001: ID_S_192fd704_45804608_E <= 8'b00010000; 4'b1010: ID_S_192fd704_45804608_E <= 8'b00001000; 4'b1011: ID_S_192fd704_45804608_E <= 8'b00000011; 4'b1100: ID_S_192fd704_45804608_E <= 8'b01000110; 4'b1101: ID_S_192fd704_45804608_E <= 8'b00100001; 4'b1110: ID_S_192fd704_45804608_E <= 8'b00000110; 4'b1111: ID_S_192fd704_45804608_E <= 8'b00001110; endcase end endmodule    module encryptor(clock, enable, in, out, reset);   input clock; input enable; input reset; input [7:0] in; output [7:0] out;             reg ID_S_2b606_61_E; reg ID_S_2b607_62_E; reg ID_S_2b608_63_E; reg ID_S_2b609_64_E; reg ID_S_2b60a_65_E; reg ID_S_2b60b_66_E; reg ID_S_2b60c_67_E; reg ID_S_2b60d_68_E; reg ID_S_2b60e_69_E; reg ID_S_2b60f_6a_E; reg ID_S_2b610_6b_E; reg ID_S_2b611_6c_E; reg ID_S_2b612_6d_E; reg ID_S_2b613_6e_E; reg ID_S_2b614_6f_E; reg ID_S_2b615_70_E; reg ID_S_2b616_71_E; reg ID_S_2b617_72_E; reg ID_S_2b618_73_E; reg ID_S_2b619_74_E; reg ID_S_2b61a_75_E; reg ID_S_2b61b_76_E; reg ID_S_2b61c_77_E; reg ID_S_2b61d_78_E; always @(posedge clock) begin ID_S_2b606_61_E <= ID_S_2b607_62_E; ID_S_2b608_63_E <= ~ID_S_2b60b_66_E; ID_S_2b60a_65_E <= ID_S_2b617_72_E << ~ID_S_2b61a_75_E; ID_S_2b609_64_E <= ID_S_2b606_61_E & ~ID_S_2b607_62_E; ID_S_2b607_62_E <= ~(ID_S_2b617_72_E | ID_S_2b619_74_E); ID_S_2b61d_78_E <= (ID_S_2b617_72_E ^ ID_S_2b60d_68_E) & (ID_S_2b617_72_E | ID_S_2b619_74_E) | ~ID_S_2b60d_68_E; ID_S_2b61b_76_E <= (ID_S_2b610_6b_E < ID_S_2b61b_76_E) ? ID_S_2b61d_78_E : ID_S_2b60a_65_E; ID_S_2b61a_75_E <= ~(ID_S_2b614_6f_E & ID_S_2b615_70_E ^ ID_S_2b60b_66_E | ~ID_S_2b616_71_E & ID_S_2b614_6f_E); ID_S_2b619_74_E <= ~(ID_S_2b60c_67_E >> ID_S_2b607_62_E); ID_S_2b617_72_E <= (ID_S_2b61a_75_E) ? ID_S_2b61a_75_E : ID_S_2b614_6f_E; ID_S_2b612_6d_E <= (ID_S_2b619_74_E & ~ID_S_2b60a_65_E); ID_S_2b60e_69_E <= ID_S_2b609_64_E & ID_S_2b61a_75_E + 1 | (ID_S_2b619_74_E & (ID_S_2b61a_75_E + 1 + (ID_S_2b606_61_E | ~ID_S_2b607_62_E - ID_S_2b608_63_E))); ID_S_2b60a_65_E <= ID_S_2b619_74_E ^ ID_S_2b60b_66_E & ID_S_2b608_63_E | ID_S_2b607_62_E & ID_S_2b613_6e_E & (ID_S_2b617_72_E | ~ID_S_2b60f_6a_E ^ ID_S_2b611_6c_E | ~ID_S_2b612_6d_E); end initial begin ID_S_2b606_61_E = 1'b0; ID_S_2b607_62_E = 1'b1; ID_S_2b608_63_E = 1'b0; ID_S_2b609_64_E = 1'b0; ID_S_2b60a_65_E = 1'b0; ID_S_2b60b_66_E = 1'b1; ID_S_2b60c_67_E = 1'b0; ID_S_2b60d_68_E = 1'b1; ID_S_2b60e_69_E = 1'b1; ID_S_2b60f_6a_E = 1'b0; ID_S_2b610_6b_E = 1'b0; ID_S_2b611_6c_E = 1'b1; ID_S_2b612_6d_E = 1'b1; ID_S_2b613_6e_E = 1'b0; ID_S_2b614_6f_E = 1'b1; ID_S_2b615_70_E = 1'b0; ID_S_2b616_71_E = 1'b0; ID_S_2b617_72_E = 1'b0; ID_S_2b618_73_E = 1'b1; ID_S_2b619_74_E = 1'b0; ID_S_2b61a_75_E = 1'b0; ID_S_2b61b_76_E = 1'b1; ID_S_2b61c_77_E = 1'b1; ID_S_2b61d_78_E = 1'b0; end wire ID_S_b885bf6_7e78880b_E; wire ID_S_b886037_7e749288_E; wire ID_S_b886478_7e709b09_E; wire ID_S_b8868b9_7e6ca78e_E; wire ID_S_b886cfa_7e68ae0f_E; wire ID_S_b88713b_7e64b48c_E; wire ID_S_b88757c_7e60bd0d_E; wire ID_S_b8879bd_7e5ccd83_E; wire ID_S_b885bf7_7e788808_E; wire ID_S_b886038_7e74928b_E; wire ID_S_b886479_7e709b0a_E; wire ID_S_b8868ba_7e6ca78d_E; wire ID_S_b886cfb_7e68ae0c_E; wire ID_S_b88713c_7e64b48f_E; wire ID_S_b88757d_7e60bd0e_E; wire ID_S_b8879be_7e5ccd80_E; wire ID_S_b885bf8_7e788809_E; wire ID_S_b886039_7e74928a_E; wire ID_S_b88647a_7e709b0b_E; wire ID_S_b8868bb_7e6ca78c_E; wire ID_S_b886cfc_7e68ae0d_E; wire ID_S_b88713d_7e64b48e_E; wire ID_S_b88757e_7e60bd0f_E; wire ID_S_b8879bf_7e5ccd81_E; wire ID_S_b885bf9_7e78880e_E; wire ID_S_b88603a_7e74928d_E; wire ID_S_b88647b_7e709b0c_E; wire ID_S_b8868bc_7e6ca78b_E; wire ID_S_b886cfd_7e68ae0a_E; wire ID_S_b88713e_7e64b489_E; wire ID_S_b88757f_7e60bd08_E; wire ID_S_b8879c0_7e5ccd86_E; wire ID_S_b885bfa_7e78880f_E; wire ID_S_b88603b_7e74928c_E; wire ID_S_b88647c_7e709b0d_E; wire ID_S_b8868bd_7e6ca78a_E; wire ID_S_b886cfe_7e68ae0b_E; wire ID_S_b88713f_7e64b488_E; wire ID_S_b887580_7e60bd09_E; wire ID_S_b8879c1_7e5ccd87_E; wire ID_S_b885bfb_7e78880c_E; wire ID_S_b88603c_7e74928f_E; wire ID_S_b88647d_7e709b0e_E; wire ID_S_b8868be_7e6ca789_E; wire ID_S_b886cff_7e68ae08_E; wire ID_S_b887140_7e64b48b_E; wire ID_S_b887581_7e60bd0a_E; wire ID_S_b8879c2_7e5ccd84_E; wire ID_S_b887dfe_7e58c402_E; wire ID_S_b88823f_7e54de81_E; wire ID_S_b888680_7e50d700_E; wire ID_S_b888ac1_7e4ceb87_E; wire ID_S_b888f02_7e48e206_E; wire ID_S_b889343_7e44f885_E; wire ID_S_b889784_7e40f104_E; wire ID_S_b889bc5_7e3c1998_E; wire ID_S_b887dff_7e58c401_E; wire ID_S_b888240_7e54de82_E; wire ID_S_b888681_7e50d703_E; wire ID_S_b888ac2_7e4ceb84_E; wire ID_S_b888f03_7e48e205_E; wire ID_S_b889344_7e44f886_E; wire ID_S_b889785_7e40f107_E; wire ID_S_b889bc6_7e3c199b_E; wire ID_S_b887e00_7e58c400_E; wire ID_S_b888241_7e54de83_E; wire ID_S_b888682_7e50d702_E; wire ID_S_b888ac3_7e4ceb85_E; wire ID_S_b888f04_7e48e204_E; wire ID_S_b889345_7e44f887_E; wire ID_S_b889786_7e40f106_E; wire ID_S_b889bc7_7e3c199a_E; wire ID_S_b887e01_7e58c407_E; wire ID_S_b888242_7e54de84_E; wire ID_S_b888683_7e50d705_E; wire ID_S_b888ac4_7e4ceb82_E; wire ID_S_b888f05_7e48e203_E; wire ID_S_b889346_7e44f880_E; wire ID_S_b889787_7e40f101_E; wire ID_S_b889bc8_7e3c199d_E; wire ID_S_b887e02_7e58c406_E; wire ID_S_b888243_7e54de85_E; wire ID_S_b888684_7e50d704_E; wire ID_S_b888ac5_7e4ceb83_E; wire ID_S_b888f06_7e48e202_E; wire ID_S_b889347_7e44f881_E; wire ID_S_b889788_7e40f100_E; wire ID_S_b889bc9_7e3c199c_E; wire ID_S_b887e03_7e58c405_E; wire ID_S_b888244_7e54de86_E; wire ID_S_b888685_7e50d707_E; wire ID_S_b888ac6_7e4ceb80_E; wire ID_S_b888f07_7e48e201_E; wire ID_S_b889348_7e44f882_E; wire ID_S_b889789_7e40f103_E; wire ID_S_b889bca_7e3c199f_E; ID_S_7efb9f9e_394c97fa_E ID_S_597927_7ffc6fbe_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b606_61_E,ID_S_2b607_62_E,ID_S_2b608_63_E,ID_S_2b609_64_E}), .ID_S_192fd704_45804608_E({ID_S_b885bf6_7e78880b_E,ID_S_b886037_7e749288_E,ID_S_b886478_7e709b09_E,ID_S_b8868b9_7e6ca78e_E,ID_S_b886cfa_7e68ae0f_E,ID_S_b88713b_7e64b48c_E,ID_S_b88757c_7e60bd0d_E,ID_S_b8879bd_7e5ccd83_E})); ID_S_7efb9f9e_394c97fa_E ID_S_597928_7ffc6fbf_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b60a_65_E,ID_S_2b60b_66_E,ID_S_2b60c_67_E,ID_S_2b60d_68_E}), .ID_S_192fd704_45804608_E({ID_S_b885bf7_7e788808_E,ID_S_b886038_7e74928b_E,ID_S_b886479_7e709b0a_E,ID_S_b8868ba_7e6ca78d_E,ID_S_b886cfb_7e68ae0c_E,ID_S_b88713c_7e64b48f_E,ID_S_b88757d_7e60bd0e_E,ID_S_b8879be_7e5ccd80_E})); ID_S_7efb9f9e_394c97fa_E ID_S_597929_7ffc6fbc_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b60e_69_E,ID_S_2b60f_6a_E,ID_S_2b610_6b_E,ID_S_2b611_6c_E}), .ID_S_192fd704_45804608_E({ID_S_b885bf8_7e788809_E,ID_S_b886039_7e74928a_E,ID_S_b88647a_7e709b0b_E,ID_S_b8868bb_7e6ca78c_E,ID_S_b886cfc_7e68ae0d_E,ID_S_b88713d_7e64b48e_E,ID_S_b88757e_7e60bd0f_E,ID_S_b8879bf_7e5ccd81_E})); ID_S_7efb9f9e_394c97fa_E ID_S_59792a_7ffc6fbd_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b612_6d_E,ID_S_2b613_6e_E,ID_S_2b614_6f_E,ID_S_2b615_70_E}), .ID_S_192fd704_45804608_E({ID_S_b885bf9_7e78880e_E,ID_S_b88603a_7e74928d_E,ID_S_b88647b_7e709b0c_E,ID_S_b8868bc_7e6ca78b_E,ID_S_b886cfd_7e68ae0a_E,ID_S_b88713e_7e64b489_E,ID_S_b88757f_7e60bd08_E,ID_S_b8879c0_7e5ccd86_E})); ID_S_7efb9f9e_394c97fa_E ID_S_59792b_7ffc6fba_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b616_71_E,ID_S_2b617_72_E,ID_S_2b618_73_E,ID_S_2b619_74_E}), .ID_S_192fd704_45804608_E({ID_S_b885bfa_7e78880f_E,ID_S_b88603b_7e74928c_E,ID_S_b88647c_7e709b0d_E,ID_S_b8868bd_7e6ca78a_E,ID_S_b886cfe_7e68ae0b_E,ID_S_b88713f_7e64b488_E,ID_S_b887580_7e60bd09_E,ID_S_b8879c1_7e5ccd87_E})); ID_S_7efb9f9e_394c97fa_E ID_S_59792c_7ffc6fbb_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b61a_75_E,ID_S_2b61b_76_E,ID_S_2b61c_77_E,ID_S_2b61d_78_E}), .ID_S_192fd704_45804608_E({ID_S_b885bfb_7e78880c_E,ID_S_b88603c_7e74928f_E,ID_S_b88647d_7e709b0e_E,ID_S_b8868be_7e6ca789_E,ID_S_b886cff_7e68ae08_E,ID_S_b887140_7e64b48b_E,ID_S_b887581_7e60bd0a_E,ID_S_b8879c2_7e5ccd84_E})); ID_S_7efb9f9e_394c97fa_E ID_S_59792d_7ffc6fb8_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b606_61_E,ID_S_2b607_62_E,ID_S_2b608_63_E,ID_S_2b609_64_E}), .ID_S_192fd704_45804608_E({ID_S_b887dfe_7e58c402_E,ID_S_b88823f_7e54de81_E,ID_S_b888680_7e50d700_E,ID_S_b888ac1_7e4ceb87_E,ID_S_b888f02_7e48e206_E,ID_S_b889343_7e44f885_E,ID_S_b889784_7e40f104_E,ID_S_b889bc5_7e3c1998_E})); ID_S_7efb9f9e_394c97fa_E ID_S_59792e_7ffc6fb9_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b60a_65_E,ID_S_2b60b_66_E,ID_S_2b60c_67_E,ID_S_2b60d_68_E}), .ID_S_192fd704_45804608_E({ID_S_b887dff_7e58c401_E,ID_S_b888240_7e54de82_E,ID_S_b888681_7e50d703_E,ID_S_b888ac2_7e4ceb84_E,ID_S_b888f03_7e48e205_E,ID_S_b889344_7e44f886_E,ID_S_b889785_7e40f107_E,ID_S_b889bc6_7e3c199b_E})); ID_S_7efb9f9e_394c97fa_E ID_S_59792f_7ffc6fb6_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b60e_69_E,ID_S_2b60f_6a_E,ID_S_2b610_6b_E,ID_S_2b611_6c_E}), .ID_S_192fd704_45804608_E({ID_S_b887e00_7e58c400_E,ID_S_b888241_7e54de83_E,ID_S_b888682_7e50d702_E,ID_S_b888ac3_7e4ceb85_E,ID_S_b888f04_7e48e204_E,ID_S_b889345_7e44f887_E,ID_S_b889786_7e40f106_E,ID_S_b889bc7_7e3c199a_E})); ID_S_7efb9f9e_394c97fa_E ID_S_597930_7ffc6fb7_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b612_6d_E,ID_S_2b613_6e_E,ID_S_2b614_6f_E,ID_S_2b615_70_E}), .ID_S_192fd704_45804608_E({ID_S_b887e01_7e58c407_E,ID_S_b888242_7e54de84_E,ID_S_b888683_7e50d705_E,ID_S_b888ac4_7e4ceb82_E,ID_S_b888f05_7e48e203_E,ID_S_b889346_7e44f880_E,ID_S_b889787_7e40f101_E,ID_S_b889bc8_7e3c199d_E})); ID_S_7efb9f9e_394c97fa_E ID_S_597938_7ffc6fcf_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b616_71_E,ID_S_2b617_72_E,ID_S_2b618_73_E,ID_S_2b619_74_E}), .ID_S_192fd704_45804608_E({ID_S_b887e02_7e58c406_E,ID_S_b888243_7e54de85_E,ID_S_b888684_7e50d704_E,ID_S_b888ac5_7e4ceb83_E,ID_S_b888f06_7e48e202_E,ID_S_b889347_7e44f881_E,ID_S_b889788_7e40f100_E,ID_S_b889bc9_7e3c199c_E})); ID_S_7efb9f9e_394c97fa_E ID_S_597939_7ffc6fcc_E (.clock(clock), .ID_S_108d5742_7edd6db7_E({ID_S_2b61a_75_E,ID_S_2b61b_76_E,ID_S_2b61c_77_E,ID_S_2b61d_78_E}), .ID_S_192fd704_45804608_E({ID_S_b887e03_7e58c405_E,ID_S_b888244_7e54de86_E,ID_S_b888685_7e50d707_E,ID_S_b888ac6_7e4ceb80_E,ID_S_b888f07_7e48e201_E,ID_S_b889348_7e44f882_E,ID_S_b889789_7e40f103_E,ID_S_b889bca_7e3c199f_E})); wire ID_S_b888d0c_7e4cf3ec_E; wire ID_S_597906_7ffc77bd_E, ID_S_597907_7ffc77bc_E, ID_S_597908_7ffc77bf_E; wire ID_S_597759_7ffcdfa8_E, ID_S_59775a_7ffcdfa9_E, ID_S_59775b_7ffcdfaa_E; wire ID_S_5977fe_7ffcb7a5_E, ID_S_5977ff_7ffcb7a4_E, ID_S_597800_7ffcb7a7_E, ID_S_597801_7ffcb7a6_E; wire ID_S_5978c4_7ffc87a3_E, ID_S_5978c5_7ffc87a2_E, ID_S_5978c6_7ffc87a1_E, ID_S_5978c7_7ffc87a0_E, ID_S_5978c8_7ffc87a7_E; wire [3:0] ID_S_302b34b2_b38ae8c_E; reg [3:0] ID_S_7c9e679b_1f355465_E; ID_S_5d0f61ec_7e71e69b_E ID_S_597882_7ffc97a1_E (.ID_S_2b616_71_E(ID_S_597906_7ffc77bd_E), .ID_S_2b609_64_E(ID_S_597759_7ffcdfa8_E), .clock(clock), .reset(reset)); ID_S_5d0f61ec_7e71e69b_E ID_S_597883_7ffc97a0_E (.ID_S_2b616_71_E(ID_S_597907_7ffc77bc_E), .ID_S_2b609_64_E(ID_S_59775a_7ffcdfa9_E), .clock(clock), .reset(reset)); ID_S_5d0f61ec_7e71e69b_E ID_S_597884_7ffc97a3_E (.ID_S_2b616_71_E(ID_S_597908_7ffc77bf_E), .ID_S_2b609_64_E(ID_S_59775b_7ffcdfaa_E), .clock(clock), .reset(reset)); initial begin ID_S_7c9e679b_1f355465_E = 4'b0110; end assign ID_S_5977fe_7ffcb7a5_E = ID_S_7c9e679b_1f355465_E[3]; assign ID_S_5977ff_7ffcb7a4_E = ID_S_7c9e679b_1f355465_E[2]; assign ID_S_597800_7ffcb7a7_E = ID_S_7c9e679b_1f355465_E[1]; assign ID_S_597801_7ffcb7a6_E = ID_S_7c9e679b_1f355465_E[0]; assign ID_S_597759_7ffcdfa8_E = ((~ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ID_S_597908_7ffc77bf_E & ~ID_S_5977fe_7ffcb7a5_E)&((ID_S_5977ff_7ffcb7a4_E&ID_S_597800_7ffcb7a7_E) | (~ID_S_597800_7ffcb7a7_E&ID_S_597801_7ffcb7a6_E) | (ID_S_597800_7ffcb7a7_E&~ID_S_597801_7ffcb7a6_E))) | ((~ID_S_597906_7ffc77bd_E & ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E & ~ID_S_5977fe_7ffcb7a5_E)&((ID_S_5977ff_7ffcb7a4_E&ID_S_597801_7ffcb7a6_E) | (ID_S_5977ff_7ffcb7a4_E&ID_S_597800_7ffcb7a7_E&~ID_S_597801_7ffcb7a6_E) | (~ID_S_5977ff_7ffcb7a4_E&~ID_S_597800_7ffcb7a7_E&ID_S_597801_7ffcb7a6_E))) | ID_S_597906_7ffc77bd_E; assign ID_S_59775a_7ffcdfa9_E = (~ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ID_S_597908_7ffc77bf_E & ~ID_S_5977fe_7ffcb7a5_E & ID_S_5977ff_7ffcb7a4_E & ~ID_S_597800_7ffcb7a7_E & ~ID_S_597801_7ffcb7a6_E) | (~ID_S_597906_7ffc77bd_E & ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E & ~(~ID_S_5977fe_7ffcb7a5_E & ~ID_S_5977ff_7ffcb7a4_E & ~ID_S_597800_7ffcb7a7_E & ID_S_597801_7ffcb7a6_E)) | (ID_S_597906_7ffc77bd_E & ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E); assign ID_S_59775b_7ffcdfaa_E = (~ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E & ~ID_S_5977fe_7ffcb7a5_E & ~ID_S_5977ff_7ffcb7a4_E & ID_S_597800_7ffcb7a7_E & ID_S_597801_7ffcb7a6_E) | (~ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ID_S_597908_7ffc77bf_E & ((~ID_S_5977fe_7ffcb7a5_E & ~ID_S_5977ff_7ffcb7a4_E & ~ID_S_597800_7ffcb7a7_E & ~ID_S_597801_7ffcb7a6_E) | (~ID_S_5977fe_7ffcb7a5_E & ~ID_S_5977ff_7ffcb7a4_E & ID_S_597800_7ffcb7a7_E & ID_S_597801_7ffcb7a6_E) | ID_S_5977fe_7ffcb7a5_E)) | (~ID_S_597906_7ffc77bd_E & ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E & ~ID_S_5977fe_7ffcb7a5_E & ~ID_S_5977ff_7ffcb7a4_E & ~ID_S_597800_7ffcb7a7_E & ID_S_597801_7ffcb7a6_E) | (ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ID_S_597908_7ffc77bf_E); assign ID_S_5978c4_7ffc87a3_E = ~ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E; assign ID_S_5978c5_7ffc87a2_E = ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E; assign ID_S_5978c6_7ffc87a1_E = (ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E & ID_S_597908_7ffc77bf_E) | (~ID_S_597906_7ffc77bd_E & ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E); assign ID_S_5978c7_7ffc87a0_E = ID_S_597906_7ffc77bd_E & ID_S_597907_7ffc77bc_E & ~ID_S_597908_7ffc77bf_E; assign ID_S_5978c8_7ffc87a7_E = (ID_S_597906_7ffc77bd_E & ~ID_S_597908_7ffc77bf_E) | (ID_S_597906_7ffc77bd_E & ~ID_S_597907_7ffc77bc_E); assign ID_S_302b34b2_b38ae8c_E = {ID_S_5978c4_7ffc87a3_E,ID_S_5978c5_7ffc87a2_E,ID_S_5978c6_7ffc87a1_E,ID_S_5978c7_7ffc87a0_E}; assign ID_S_b888d0c_7e4cf3ec_E = ID_S_5978c8_7ffc87a7_E;         reg [7:0] ID_S_5976e8_7ffd07c6_E;   reg [7:0] ID_S_5976ef_7ffd07c9_E;     always @(posedge clock or posedge reset) begin     if (reset) begin ID_S_5976e8_7ffd07c6_E <= 8'b00000000; ID_S_5976ef_7ffd07c9_E <= 8'b01101001;   end   else if (enable) begin ID_S_5976e8_7ffd07c6_E <= (in ^ ID_S_5976ef_7ffd07c9_E);   ID_S_5976ef_7ffd07c9_E <= (ID_S_5976ef_7ffd07c9_E - 2);   end end   assign out = ID_S_5976e8_7ffd07c6_E + (     ({ID_S_7c9e679b_1f355465_E, ID_S_302b34b2_b38ae8c_E} - {ID_S_7c9e679b_1f355465_E, ID_S_302b34b2_b38ae8c_E}) + ({ID_S_b885bf6_7e78880b_E,ID_S_b886037_7e749288_E,ID_S_b886478_7e709b09_E,ID_S_b8868b9_7e6ca78e_E,ID_S_b886cfa_7e68ae0f_E,ID_S_b88713b_7e64b48c_E,ID_S_b88757c_7e60bd0d_E,ID_S_b8879bd_7e5ccd83_E} - {ID_S_b885bf6_7e78880b_E,ID_S_b886037_7e749288_E,ID_S_b886478_7e709b09_E,ID_S_b8868b9_7e6ca78e_E,ID_S_b886cfa_7e68ae0f_E,ID_S_b88713b_7e64b48c_E,ID_S_b88757c_7e60bd0d_E,ID_S_b8879bd_7e5ccd83_E}) + ({ID_S_b885bf7_7e788808_E,ID_S_b886038_7e74928b_E,ID_S_b886479_7e709b0a_E,ID_S_b8868ba_7e6ca78d_E,ID_S_b886cfb_7e68ae0c_E,ID_S_b88713c_7e64b48f_E,ID_S_b88757d_7e60bd0e_E,ID_S_b8879be_7e5ccd80_E} - {ID_S_b885bf7_7e788808_E,ID_S_b886038_7e74928b_E,ID_S_b886479_7e709b0a_E,ID_S_b8868ba_7e6ca78d_E,ID_S_b886cfb_7e68ae0c_E,ID_S_b88713c_7e64b48f_E,ID_S_b88757d_7e60bd0e_E,ID_S_b8879be_7e5ccd80_E}) + ({ID_S_b885bf8_7e788809_E,ID_S_b886039_7e74928a_E,ID_S_b88647a_7e709b0b_E,ID_S_b8868bb_7e6ca78c_E,ID_S_b886cfc_7e68ae0d_E,ID_S_b88713d_7e64b48e_E,ID_S_b88757e_7e60bd0f_E,ID_S_b8879bf_7e5ccd81_E} - {ID_S_b885bf8_7e788809_E,ID_S_b886039_7e74928a_E,ID_S_b88647a_7e709b0b_E,ID_S_b8868bb_7e6ca78c_E,ID_S_b886cfc_7e68ae0d_E,ID_S_b88713d_7e64b48e_E,ID_S_b88757e_7e60bd0f_E,ID_S_b8879bf_7e5ccd81_E}) + ({ID_S_b885bf9_7e78880e_E,ID_S_b88603a_7e74928d_E,ID_S_b88647b_7e709b0c_E,ID_S_b8868bc_7e6ca78b_E,ID_S_b886cfd_7e68ae0a_E,ID_S_b88713e_7e64b489_E,ID_S_b88757f_7e60bd08_E,ID_S_b8879c0_7e5ccd86_E} - {ID_S_b885bf9_7e78880e_E,ID_S_b88603a_7e74928d_E,ID_S_b88647b_7e709b0c_E,ID_S_b8868bc_7e6ca78b_E,ID_S_b886cfd_7e68ae0a_E,ID_S_b88713e_7e64b489_E,ID_S_b88757f_7e60bd08_E,ID_S_b8879c0_7e5ccd86_E}) + ({ID_S_b885bfa_7e78880f_E,ID_S_b88603b_7e74928c_E,ID_S_b88647c_7e709b0d_E,ID_S_b8868bd_7e6ca78a_E,ID_S_b886cfe_7e68ae0b_E,ID_S_b88713f_7e64b488_E,ID_S_b887580_7e60bd09_E,ID_S_b8879c1_7e5ccd87_E} - {ID_S_b885bfa_7e78880f_E,ID_S_b88603b_7e74928c_E,ID_S_b88647c_7e709b0d_E,ID_S_b8868bd_7e6ca78a_E,ID_S_b886cfe_7e68ae0b_E,ID_S_b88713f_7e64b488_E,ID_S_b887580_7e60bd09_E,ID_S_b8879c1_7e5ccd87_E}) + ({ID_S_b885bfb_7e78880c_E,ID_S_b88603c_7e74928f_E,ID_S_b88647d_7e709b0e_E,ID_S_b8868be_7e6ca789_E,ID_S_b886cff_7e68ae08_E,ID_S_b887140_7e64b48b_E,ID_S_b887581_7e60bd0a_E,ID_S_b8879c2_7e5ccd84_E} - {ID_S_b885bfb_7e78880c_E,ID_S_b88603c_7e74928f_E,ID_S_b88647d_7e709b0e_E,ID_S_b8868be_7e6ca789_E,ID_S_b886cff_7e68ae08_E,ID_S_b887140_7e64b48b_E,ID_S_b887581_7e60bd0a_E,ID_S_b8879c2_7e5ccd84_E}) + ({ID_S_b887dfe_7e58c402_E,ID_S_b88823f_7e54de81_E,ID_S_b888680_7e50d700_E,ID_S_b888ac1_7e4ceb87_E,ID_S_b888f02_7e48e206_E,ID_S_b889343_7e44f885_E,ID_S_b889784_7e40f104_E,ID_S_b889bc5_7e3c1998_E} - {ID_S_b887dfe_7e58c402_E,ID_S_b88823f_7e54de81_E,ID_S_b888680_7e50d700_E,ID_S_b888ac1_7e4ceb87_E,ID_S_b888f02_7e48e206_E,ID_S_b889343_7e44f885_E,ID_S_b889784_7e40f104_E,ID_S_b889bc5_7e3c1998_E}) + ({ID_S_b887dff_7e58c401_E,ID_S_b888240_7e54de82_E,ID_S_b888681_7e50d703_E,ID_S_b888ac2_7e4ceb84_E,ID_S_b888f03_7e48e205_E,ID_S_b889344_7e44f886_E,ID_S_b889785_7e40f107_E,ID_S_b889bc6_7e3c199b_E} - {ID_S_b887dff_7e58c401_E,ID_S_b888240_7e54de82_E,ID_S_b888681_7e50d703_E,ID_S_b888ac2_7e4ceb84_E,ID_S_b888f03_7e48e205_E,ID_S_b889344_7e44f886_E,ID_S_b889785_7e40f107_E,ID_S_b889bc6_7e3c199b_E}) + ({ID_S_b887e00_7e58c400_E,ID_S_b888241_7e54de83_E,ID_S_b888682_7e50d702_E,ID_S_b888ac3_7e4ceb85_E,ID_S_b888f04_7e48e204_E,ID_S_b889345_7e44f887_E,ID_S_b889786_7e40f106_E,ID_S_b889bc7_7e3c199a_E} - {ID_S_b887e00_7e58c400_E,ID_S_b888241_7e54de83_E,ID_S_b888682_7e50d702_E,ID_S_b888ac3_7e4ceb85_E,ID_S_b888f04_7e48e204_E,ID_S_b889345_7e44f887_E,ID_S_b889786_7e40f106_E,ID_S_b889bc7_7e3c199a_E}) + ({ID_S_b887e01_7e58c407_E,ID_S_b888242_7e54de84_E,ID_S_b888683_7e50d705_E,ID_S_b888ac4_7e4ceb82_E,ID_S_b888f05_7e48e203_E,ID_S_b889346_7e44f880_E,ID_S_b889787_7e40f101_E,ID_S_b889bc8_7e3c199d_E} - {ID_S_b887e01_7e58c407_E,ID_S_b888242_7e54de84_E,ID_S_b888683_7e50d705_E,ID_S_b888ac4_7e4ceb82_E,ID_S_b888f05_7e48e203_E,ID_S_b889346_7e44f880_E,ID_S_b889787_7e40f101_E,ID_S_b889bc8_7e3c199d_E}) + ({ID_S_b887e02_7e58c406_E,ID_S_b888243_7e54de85_E,ID_S_b888684_7e50d704_E,ID_S_b888ac5_7e4ceb83_E,ID_S_b888f06_7e48e202_E,ID_S_b889347_7e44f881_E,ID_S_b889788_7e40f100_E,ID_S_b889bc9_7e3c199c_E} - {ID_S_b887e02_7e58c406_E,ID_S_b888243_7e54de85_E,ID_S_b888684_7e50d704_E,ID_S_b888ac5_7e4ceb83_E,ID_S_b888f06_7e48e202_E,ID_S_b889347_7e44f881_E,ID_S_b889788_7e40f100_E,ID_S_b889bc9_7e3c199c_E}) + ({ID_S_b887e03_7e58c405_E,ID_S_b888244_7e54de86_E,ID_S_b888685_7e50d707_E,ID_S_b888ac6_7e4ceb80_E,ID_S_b888f07_7e48e201_E,ID_S_b889348_7e44f882_E,ID_S_b889789_7e40f103_E,ID_S_b889bca_7e3c199f_E} - {ID_S_b887e03_7e58c405_E,ID_S_b888244_7e54de86_E,ID_S_b888685_7e50d707_E,ID_S_b888ac6_7e4ceb80_E,ID_S_b888f07_7e48e201_E,ID_S_b889348_7e44f882_E,ID_S_b889789_7e40f103_E,ID_S_b889bca_7e3c199f_E}) ); endmodule 